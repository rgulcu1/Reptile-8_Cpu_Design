module ControlUnit(opcode,clk,Armux,MemLoad,PcLoad,PcInc,RegLoad,ZfLoad,mux,IrLoad);

endmodule
